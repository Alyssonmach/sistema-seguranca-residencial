// modulo de uma and de 3 entradas
module and_3entradas
(
	input A,B,C,
	output S1
);

 assign S1 = A & B & C;
 
endmodule 
// sistema de segurança residencial
// alysson machado e matheus victor