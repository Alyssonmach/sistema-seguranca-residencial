// modulo de uma or de 6 entradas
module or_6entradas
(
	input A,B,C,D,E,F,
	output S2

);

	assign S2 = A | B | C | D | E | F; 


endmodule 
// sistema de segurança residencial
// alysson machado e matheus victor